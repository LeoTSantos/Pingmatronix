library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package SSDefinitions is
	type SSD_ARRAY is array (natural range<>) of std_logic_vector(0 to 6);

end package;