
package PongDefinitions is

    
    constant MAX_RACKET_Y: NATURAL := 44;
    constant MIN_RACKET_Y: NATURAL := 3;
    constant MAX_PONTOS: NATURAL := 10;

    
end package;