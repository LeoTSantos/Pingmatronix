library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.math_real.all;

package VgaDefinitions is
	constant VGA_MAX_HORIZONTAL:natural := 63;
	constant VGA_MAX_VERTICAL:natural := 47;
end package;